module MemWb(
    input  wire        clk,
    input  wire        rst,
    input  wire [9:0]  mem_control_sig,
    input  wire [31:0] mem_memval,
    input  wire [31:0] mem_alu,
    input  wire [4:0]  mem_rd,

    output reg  [9:0]  wb_control_sig,
    output reg  [31:0] wb_memval,
    output reg  [31:0] wb_alu,
    output reg  [4:0]  wb_rd
);

    always @(posedge clk or posedge rst) 
	begin
        if (rst) 
		begin
            	wb_control_sig <= 10'b0;
            	wb_memval      <= 32'b0;
            	wb_alu         <= 32'b0;
            	wb_rd          <= 5'b0;
        	end
        else 
		begin
            	wb_control_sig <= mem_control_sig;
            	wb_memval      <= mem_memval;
            	wb_alu         <= mem_alu;
            	wb_rd          <= mem_rd;
        	end
    	end

endmodule
